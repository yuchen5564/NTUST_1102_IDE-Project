* Project05: L08-P13.sp

r1 0 a 10

l1 a 0 10m ic=1

.tran 0.1ms 10ms uic

.end
