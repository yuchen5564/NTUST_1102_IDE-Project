* Project05; L07-P15.sp

v1 a 0 dc 10

vdr1 c 0 dc 0

r1 a b 1k

c1 b c 1u ic=0

.tran 0.1ms 10ms uic

.end

