* Project05: L07-P17.sp

vdr1 0 b dc 0

r1 b a 1k

c1 a 0 1u ic=10

.tran 0.1ms 10ms uic

.end
