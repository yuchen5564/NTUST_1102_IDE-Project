* Project05: L08-P11.sp

v1 a 0 dc 10

r1 a b 10

l1 b 0 10m ic=0

.tran 0.1ms 10ms uic

.end
